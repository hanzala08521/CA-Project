`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/25/2024 01:33:54 PM
// Design Name: 
// Module Name: ImmGen
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ImmGen
(
    input [31:0] instruc,
    output reg [63:0] imm_data
);

wire [6:0] opcode;
assign opcode = instruc[6:0];
reg [63:0] imm_data_reg;

always @(*)
begin
    case (opcode)
        7'b0000011: imm_data =  {{52{instruc[31]}}, instruc [31:20]}; //I
        7'b0100011: imm_data = {{52{instruc[31]}}, instruc [31:25], instruc [11:7]}; //S
        7'b1100011: imm_data = {{52{instruc[31]}}, instruc [31] , instruc [7], instruc [30:25], instruc [11:8]};
        7'b0010011: imm_data = {    {52{instruc[31]}}, instruc[31:20] };
        default : imm_data = 64'd0;
    endcase
end

endmodule